library verilog;
use verilog.vl_types.all;
entity RCA_tb is
end RCA_tb;
