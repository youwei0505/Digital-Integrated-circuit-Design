module FA(s, c_out, x, y, c_in);
input x, y, c_in;
output s, c_out;
wire s1, c1, c2;

/*
	Write Your Design Here ~
*/

//By Order
HA HA1(s1,c1,x,y);
HA HA2(s,c2,c_in,s1);
or or1(c_out,c2,c1);

endmodule

